module top (
	input clk,
	input key,
	output [7:0] led
);
    assign led = 8'b11111111;
    



endmodule
